module ex();
  
  
endmodule