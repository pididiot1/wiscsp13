/* $Author: karu $ */
/* $LastChangedDate: 2009-03-04 23:09:45 -0600 (Wed, 04 Mar 2009) $ */
/* $Rev: 45 $ */
module proc (/*AUTOARG*/
   // Outputs
   err, 
   // Inputs
   clk, rst
   );

   input clk;
   input rst;

   output err;

   // None of the above lines can be modified

   // OR all the err ouputs for every sub-module and assign it as this
   // err output
   
   // As desribed in the homeworks, use the err signal to trap corner
   // cases that you think are illegal in your statemachines
   
   
   /* your code here */
   infetch fetch(
                  //Inputs
                  .clk(clk), .rst(rst)
                  //Outputs
                  );
   id decode(
                  //Inputs
                  .clk(clk), .rst(rst)
                  //Outputs
                  );
   ex execute(
                  //Inputs
                  //Outputs
                  );
   mem memfetch(
                  //Inputs
                  .clk(clk), .rst(rst)
                  //Outputs
                  );
   wb writeback(
                  //Inputs
                  //Outputs
                  );
   
endmodule // proc
// DUMMY LINE FOR REV CONTROL :0: