module wb();
  
  
endmodule