module claAdder(Sum, G, P, Cout, Cprev, A, B, Cin);

output [15:0] Sum, G, P;
output Cout, Cprev;
input [15:0] A, B;
input Cin;

wire c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15;

assign P[0] = A[0] | B[0];
assign G[0] = A[0] & B[0];
assign P[1] = A[1] | B[1];
assign G[1] = A[1] & B[1];
assign P[2] = A[2] | B[2];
assign G[2] = A[2] & B[2];
assign P[3] = A[3] | B[3];
assign G[3] = A[3] & B[3];
assign P[4] = A[4] | B[4];
assign G[4] = A[4] & B[4];
assign P[5] = A[5] | B[5];
assign G[5] = A[5] & B[5];
assign P[6] = A[6] | B[6];
assign G[6] = A[6] & B[6];
assign P[7] = A[7] | B[7];
assign G[7] = A[7] & B[7];
assign P[8] = A[8] | B[8];
assign G[8] = A[8] & B[8];
assign P[9] = A[9] | B[9];
assign G[9] = A[9] & B[9];
assign P[10] = A[10] | B[10];
assign G[10] = A[10] & B[10];
assign P[11] = A[11] | B[11];
assign G[11] = A[11] & B[11];
assign P[12] = A[12] | B[12];
assign G[12] = A[12] & B[12];
assign P[13] = A[13] | B[13];
assign G[13] = A[13] & B[13];
assign P[14] = A[14] | B[14];
assign G[14] = A[14] & B[14];
assign P[15] = A[15] | B[15];
assign G[15] = A[15] & B[15];

assign c1 = G[0] | (P[0] & Cin);
assign c2 = G[1] | (P[1] & G[0]) | (P[1] & P[0] & Cin);
assign c3 = G[2]| (P[2] & G[1]) | (P[2] & P[1] & G[0]) | (P[2] & P[1] & P[0] & Cin);
assign c4 = G[3]| (P[3] & G[2]) | (P[3] & P[2] & G[1]) | (P[3] & P[2] & P[1] & G[0]) | (P[3] & P[2] & P[1] & P[0] & Cin);
assign c5 = G[4] | (P[4] & G[3]) | (P[4] & P[3] & G[2]) | (P[4] & P[3] & P[2] & G[1]) | (P[4] & P[3] & P[2] & P[1] & G[0]) | (P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c6 = G[5] | (P[5] & G[4]) | (P[5] & P[4] & G[3]) | (P[5] & P[4] & P[3] & G[2]) | (P[5] & P[4] & P[3] & P[2] & G[1]) | (P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c7 = G[6] | (P[6] & G[5]) | (P[6] & P[5] & G[4]) | (P[6] & P[5] & P[4] & G[3]) | (P[6] & P[5] & P[4] & P[3] & G[2]) | (P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c8 = G[7] | (P[7] & G[6]) | (P[7] & P[6] & G[5]) | (P[7] & P[6] & P[5] & G[4]) | (P[7] & P[6] & P[5] & P[4] & G[3]) | (P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c9 = G[8] | (P[8] & G[7]) | (P[8] & P[7] & G[6]) | (P[8] & P[7] & P[6] & G[5]) | (P[8] & P[7] & P[6] & P[5] & G[4]) | (P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c10 = G[9] | (P[9] & G[8]) | (P[9] & P[8] & G[7]) | (P[9] & P[8] & P[7] & G[6]) | (P[9] & P[8] & P[7] & P[6] & G[5]) | (P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c11 = G[10] | (P[10] & G[9]) | (P[10] & P[9] & G[8]) | (P[10] & P[9] & P[8] & G[7]) | (P[10] & P[9] & P[8] & P[7] & G[6]) | (P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c12 = G[11] | (P[11] & G[10]) | (P[11] & P[10] & G[9]) | (P[11] & P[10] & P[9] & G[8]) | (P[11] & P[10] & P[9] & P[8] & G[7]) | (P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c13 = G[12] | (P[12] & G[11]) | (P[12] & P[11] & G[10]) | (P[12] & P[11] & P[10] & G[9]) | (P[12] & P[11] & P[10] & P[9] & G[8]) | (P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c14 = G[13] | (P[13] & G[12]) | (P[13] & P[12] & G[11]) | (P[13] & P[12] & P[11] & G[10]) | (P[13] & P[12] & P[11] & P[10] & G[9]) | (P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign c15 = G[14] | (P[14] & G[13]) | (P[14] & P[13] & G[12]) | (P[14] & P[13] & P[12] & G[11]) | (P[14] & P[13] & P[12] & P[11] & G[10]) | (P[14] & P[13] & P[12] & P[11] & P[10] & G[9]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);
assign Cout = G[15] | (P[15] & G[14]) | (P[15] & P[14] & G[13]) | (P[15] & P[14] & P[13] & G[12]) | (P[15] & P[14] & P[13] & P[12] & G[11]) | (P[15] & P[14] & P[13] & P[12] & P[11] & G[10]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & Cin);

assign Cprev = c15;

sum zero(.sum(Sum[0]), .a(A[0]), .b(B[0]), .cin(Cin));
sum one(.sum(Sum[1]), .a(A[1]), .b(B[1]), .cin(c1));
sum two(.sum(Sum[2]), .a(A[2]), .b(B[2]), .cin(c2));
sum three(.sum(Sum[3]), .a(A[3]), .b(B[3]), .cin(c3));
sum four(.sum(Sum[4]), .a(A[4]), .b(B[4]), .cin(c4));
sum five(.sum(Sum[5]), .a(A[5]), .b(B[5]), .cin(c5));
sum six(.sum(Sum[6]), .a(A[6]), .b(B[6]), .cin(c6));
sum seven(.sum(Sum[7]), .a(A[7]), .b(B[7]), .cin(c7));
sum eight(.sum(Sum[8]), .a(A[8]), .b(B[8]), .cin(c8));
sum nine(.sum(Sum[9]), .a(A[9]), .b(B[9]), .cin(c9));
sum ten(.sum(Sum[10]), .a(A[10]), .b(B[10]), .cin(c10));
sum eleven(.sum(Sum[11]), .a(A[11]), .b(B[11]), .cin(c11));
sum twelve(.sum(Sum[12]), .a(A[12]), .b(B[12]), .cin(c12));
sum thirteen(.sum(Sum[13]), .a(A[13]), .b(B[13]), .cin(c13));
sum fourteen(.sum(Sum[14]), .a(A[14]), .b(B[14]), .cin(c14));
sum fifteen(.sum(Sum[15]), .a(A[15]), .b(B[15]), .cin(c15));

endmodule